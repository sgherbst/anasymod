`timescale 1ns/1ps

`include "svreal.sv"
//`include "math.sv"
`include "msdsl.sv"

`default_nettype none

module sim_ctrl (
    //input `DATA_TYPE_REAL(`LONG_WIDTH_REAL) primpf
);

//`PROBE_ANALOG_CTRL(primpf, top.tb_i.v_out);

//`PROBE_DIGITAL(primpf, `LONG_WIDTH_REAL);

//`PRINT_FORMAT_REAL(top.tb_i.v_out);


endmodule

`default_nettype wire